* C:\Users\mox\Desktop\Versuch2\Schematic1.sch

* Schematics Version 9.1 - Web Update 1
* Wed Oct 30 14:08:13 2013



** Analysis setup **
.tran 0.1s 2s 0 0.01s
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic1.net"
.INC "Schematic1.als"


.probe


.END
